# Language: Swedish (CP850)
# Translation by Martin Strömberg <ams@ludd.luth.se>
0.0:Väntar tills användaren trycker på en tangent från en lista av val
0.1:val
0.2:text
0.3:Specificerar vilka tangenter som är giltiga. Default är:
0.4:Visa inte valen efter prompten
0.5:Versaler skilda från gemener
0.6:**Ignorerad, för kompatibiltet med MS-DOS
0.7:Texten som ska visas som prompt
0.8:Ljud en signal när prompten visas
3.0:jn
